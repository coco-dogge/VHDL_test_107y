module cmd_rom(
	input [15:0] address,
	output [7:0] data_out,
	output DC_data
);
reg [7:0]romA[84:0];
reg [84:0]romB;
assign data_out = romA[address];
assign DC_data = romB[address];

initial
begin
		romA[0]   	<= 8'h11;
		romA[1]   	<= 8'hb1;
		romA[2]   	<= 8'h05;
		romA[3]   	<= 8'h3c;
		romA[4]   	<= 8'h3c;
		romA[5]   	<= 8'hb2;
		romA[6]   	<= 8'h05;
		romA[7]   	<= 8'h3c;
		romA[8]   	<= 8'h3c;
		romA[9]   	<= 8'hb3;
		romA[10]   	<= 8'h05;
		romA[11]   	<= 8'h3c;
		romA[12]   	<= 8'h3c;
		romA[13]   	<= 8'h05;
		romA[14]   	<= 8'h3c;
		romA[15]   	<= 8'h3c;
		romA[16]   	<= 8'hb4;
		romA[17]   	<= 8'h03;
		romA[18]   	<= 8'hc0;
		romA[19]   	<= 8'h28;
		romA[20]   	<= 8'h08;
		romA[21]   	<= 8'h04;
		romA[22]   	<= 8'hc1;
		romA[23]   	<= 8'hc0;
		romA[24]   	<= 8'hc2;
		romA[25]   	<= 8'h0d;
		romA[26]   	<= 8'h00;
		romA[27]   	<= 8'hc3;
		romA[28]   	<= 8'h8d;
		romA[29]   	<= 8'h2a;
		romA[30]   	<= 8'hc4;
		romA[31]   	<= 8'h8d;
		romA[32]   	<= 8'hee;
		romA[33]   	<= 8'hc5;
		romA[34]   	<= 8'h1a;
		romA[35]   	<= 8'h36;
		romA[36]   	<= 8'hc0;
		romA[37]   	<= 8'he0;
		romA[38]   	<= 8'h04;
		romA[39]   	<= 8'h22;
		romA[40]   	<= 8'h07;
		romA[41]   	<= 8'h0a;
		romA[42]   	<= 8'h2e;
		romA[43]   	<= 8'h30;
		romA[44]   	<= 8'h25;
		romA[45]   	<= 8'h2a;
		romA[46]   	<= 8'h28;
		romA[47]   	<= 8'h26;
		romA[48]   	<= 8'h2e;
		romA[49]   	<= 8'h3a;
		romA[50]   	<= 8'h00;
		romA[51]   	<= 8'h01;
		romA[52]   	<= 8'h03;
		romA[53]   	<= 8'h13;
		romA[54]   	<= 8'he1;
		romA[55]   	<= 8'h04;
		romA[56]   	<= 8'h16;
		romA[57]   	<= 8'h06;
		romA[58]   	<= 8'h0d;
		romA[59]   	<= 8'h2d;
		romA[60]   	<= 8'h26;
		romA[61]   	<= 8'h23;
		romA[62]   	<= 8'h27;
		romA[63]   	<= 8'h27;
		romA[64]   	<= 8'h25;
		romA[65]   	<= 8'h2d;
		romA[66]   	<= 8'h3b;
		romA[67]   	<= 8'h00;
		romA[68]   	<= 8'h01;
		romA[69]   	<= 8'h04;
		romA[70]   	<= 8'h13;
		romA[71]   	<= 8'h3a;
		romA[72]   	<= 8'h05;
		romA[73]   	<= 8'h29;
		romA[74]   	<= 8'h2a;
		romA[75]   	<= 8'h00;
		romA[76]   	<= 8'h02;	//x1	2 		0x02
		romA[77]   	<= 8'h00;
		romA[78]   	<= 8'h81;	//x2	129	0x81
		romA[79]   	<= 8'h2b;
		romA[80]   	<= 8'h00;
		romA[81]   	<= 8'h01;	//y1	1		0x01
		romA[82]   	<= 8'h00;
		romA[83]   	<= 8'ha0;	//y2	160	0xa0
		romA[84]   	<= 8'h2c;
end

initial
begin
		romB[0]   	<= 1'b0;
		romB[1]   	<= 1'b0;
		romB[2]   	<= 1'b1;
		romB[3]   	<= 1'b1;
		romB[4]   	<= 1'b1;
		romB[5]   	<= 1'b0;
		romB[6]   	<= 1'b1;
		romB[7]   	<= 1'b1;
		romB[8]   	<= 1'b1;
		romB[9]   	<= 1'b0;
		romB[10]   	<= 1'b1;
		romB[11]   	<= 1'b1;
		romB[12]   	<= 1'b1;
		romB[13]   	<= 1'b1;
		romB[14]   	<= 1'b1;
		romB[15]   	<= 1'b1;
		romB[16]   	<= 1'b0;
		romB[17]   	<= 1'b1;
		romB[18]   	<= 1'b0;
		romB[19]   	<= 1'b1;
		romB[20]   	<= 1'b1;
		romB[21]   	<= 1'b1;
		romB[22]   	<= 1'b0;
		romB[23]   	<= 1'b1;
		romB[24]   	<= 1'b0;
		romB[25]   	<= 1'b1;
		romB[26]   	<= 1'b1;
		romB[27]   	<= 1'b0;
		romB[28]   	<= 1'b1;
		romB[29]   	<= 1'b1;
		romB[30]   	<= 1'b0;
		romB[31]   	<= 1'b1;
		romB[32]   	<= 1'b1;
		romB[33]   	<= 1'b0;
		romB[34]   	<= 1'b1;
		romB[35]   	<= 1'b0;
		romB[36]   	<= 1'b1;
		romB[37]   	<= 1'b0;
		romB[38]   	<= 1'b1;
		romB[39]   	<= 1'b1;
		romB[40]   	<= 1'b1;
		romB[41]   	<= 1'b1;
		romB[42]   	<= 1'b1;
		romB[43]   	<= 1'b1;
		romB[44]   	<= 1'b1;
		romB[45]   	<= 1'b1;
		romB[46]   	<= 1'b1;
		romB[47]   	<= 1'b1;
		romB[48]   	<= 1'b1;
		romB[49]   	<= 1'b1;
		romB[50]   	<= 1'b1;
		romB[51]   	<= 1'b1;
		romB[52]   	<= 1'b1;
		romB[53]   	<= 1'b1;
		romB[54]   	<= 1'b0;
		romB[55]   	<= 1'b1;
		romB[56]   	<= 1'b1;
		romB[57]   	<= 1'b1;
		romB[58]   	<= 1'b1;
		romB[59]   	<= 1'b1;
		romB[60]   	<= 1'b1;
		romB[61]   	<= 1'b1;
		romB[62]   	<= 1'b1;
		romB[63]   	<= 1'b1;
		romB[64]   	<= 1'b1;
		romB[65]   	<= 1'b1;
		romB[66]   	<= 1'b1;
		romB[67]   	<= 1'b1;
		romB[68]   	<= 1'b1;
		romB[69]   	<= 1'b1;
		romB[70]   	<= 1'b1;
		romB[71]   	<= 1'b0;
		romB[72]   	<= 1'b1;
		romB[73]   	<= 1'b0;
		romB[74]   	<= 1'h0;
		romB[75]   	<= 1'h1;
		romB[76]   	<= 1'h1;
		romB[77]   	<= 1'h1;
		romB[78]   	<= 1'h1;
		romB[79]   	<= 1'h0;
		romB[80]   	<= 1'h1;
		romB[81]   	<= 1'h1;
		romB[82]   	<= 1'h1;
		romB[83]   	<= 1'h1;
		romB[84]   	<= 1'h0;
end

endmodule
